
module shift_reg #(
parameter delay_cycle = 1,
parameter data_width = 32
) (
	input 					clk,
	input 					rst_n,
	input [0:0] 			shin_valid_i,
	input [data_width-1:0] 	shin_data_i,
	output [0:0] 			sho_valid_o,
	output [data_width-1:0] sho_data_o
);
	reg[0:0]			buf_valid_r[delay_cycle];
	reg[data_width-1:0] buf[delay_cycle];

genvar i;
generate
for(i=0; i<delay_cycle-1; i=i+1) begin
	always @(posedge clk or negedge rst_n) begin
		if(!rst_n) begin
			buf_valid_r[i] <= 1'b1;
		end
		else if(shin_valid_i) begin
			buf_valid_r[0] <= 1'b1;
			buf[0] <= shin_data_i;
		end
		buf_valid_r[i+1] <= buf_valid_r[i];
		buf[i+1] <= buf[i];
	end
end
endgenerate

	assign sho_valid_o = buf_valid_r[delay_cycle-1];
	assign sho_data_o  = buf[delay_cycle-1];
endmodule




module shift_regs(
	input 							 clk,
	input 							 rst_n,
	input  [0:0] 					 shin_valid_i,
	input  [`SARRAY_LOAD_WIDTH-1:0]  shin_data_i,
	output [`SARRAY_H-1:0] 			 sho_valid_o,
	output [`SARRAY_LOAD_WIDTH-1:0]  sho_data_o
);



    // -------- shift_reg0

    wire [0:0]                                   s0_shin_valid_i;
    wire [`SARRAY_LOAD_WIDTH/`SARRAY_H-1:0]      s0_shin_data_i;
    wire [0:0]                                   s0_sho_valid_o;
    wire [`SARRAY_LOAD_WIDTH/`SARRAY_H-1:0]      s0_sho_data_o;

    shift_reg #(1) u_shift_reg0 (
        .clk           (clk),
        .rst_n         (rst_n),
        .shin_valid_i  (s0_shin_valid_i),
        .shin_data_i   (s0_shin_data_i),
        .sho_valid_o   (s0_sho_valid_o),
        .sho_data_o    (s0_sho_data_o)
    );

    assign s0_shin_valid_i = shin_valid_i;
    assign s0_shin_data_i = shin_data_i[(`SARRAY_LOAD_WIDTH/`SARRAY_H*1)-1:(`SARRAY_LOAD_WIDTH/`SARRAY_H*0)];
    assign sho_valid_o[0] = s0_sho_valid_o;
    assign sho_data_o[(`SARRAY_LOAD_WIDTH/`SARRAY_H*1)-1:(`SARRAY_LOAD_WIDTH/`SARRAY_H*0)] = s0_sho_data_o;



    // -------- shift_reg1

    wire [0:0]                                   s1_shin_valid_i;
    wire [`SARRAY_LOAD_WIDTH/`SARRAY_H-1:0]      s1_shin_data_i;
    wire [0:0]                                   s1_sho_valid_o;
    wire [`SARRAY_LOAD_WIDTH/`SARRAY_H-1:0]      s1_sho_data_o;

    shift_reg #(2) u_shift_reg1 (
        .clk           (clk),
        .rst_n         (rst_n),
        .shin_valid_i  (s1_shin_valid_i),
        .shin_data_i   (s1_shin_data_i),
        .sho_valid_o   (s1_sho_valid_o),
        .sho_data_o    (s1_sho_data_o)
    );

    assign s1_shin_valid_i = shin_valid_i;
    assign s1_shin_data_i = shin_data_i[(`SARRAY_LOAD_WIDTH/`SARRAY_H*2)-1:(`SARRAY_LOAD_WIDTH/`SARRAY_H*1)];
    assign sho_valid_o[1] = s1_sho_valid_o;
    assign sho_data_o[(`SARRAY_LOAD_WIDTH/`SARRAY_H*2)-1:(`SARRAY_LOAD_WIDTH/`SARRAY_H*1)] = s1_sho_data_o;



    // -------- shift_reg2

    wire [0:0]                                   s2_shin_valid_i;
    wire [`SARRAY_LOAD_WIDTH/`SARRAY_H-1:0]      s2_shin_data_i;
    wire [0:0]                                   s2_sho_valid_o;
    wire [`SARRAY_LOAD_WIDTH/`SARRAY_H-1:0]      s2_sho_data_o;

    shift_reg #(3) u_shift_reg2 (
        .clk           (clk),
        .rst_n         (rst_n),
        .shin_valid_i  (s2_shin_valid_i),
        .shin_data_i   (s2_shin_data_i),
        .sho_valid_o   (s2_sho_valid_o),
        .sho_data_o    (s2_sho_data_o)
    );

    assign s2_shin_valid_i = shin_valid_i;
    assign s2_shin_data_i = shin_data_i[(`SARRAY_LOAD_WIDTH/`SARRAY_H*3)-1:(`SARRAY_LOAD_WIDTH/`SARRAY_H*2)];
    assign sho_valid_o[2] = s2_sho_valid_o;
    assign sho_data_o[(`SARRAY_LOAD_WIDTH/`SARRAY_H*3)-1:(`SARRAY_LOAD_WIDTH/`SARRAY_H*2)] = s2_sho_data_o;



    // -------- shift_reg3

    wire [0:0]                                   s3_shin_valid_i;
    wire [`SARRAY_LOAD_WIDTH/`SARRAY_H-1:0]      s3_shin_data_i;
    wire [0:0]                                   s3_sho_valid_o;
    wire [`SARRAY_LOAD_WIDTH/`SARRAY_H-1:0]      s3_sho_data_o;

    shift_reg #(4) u_shift_reg3 (
        .clk           (clk),
        .rst_n         (rst_n),
        .shin_valid_i  (s3_shin_valid_i),
        .shin_data_i   (s3_shin_data_i),
        .sho_valid_o   (s3_sho_valid_o),
        .sho_data_o    (s3_sho_data_o)
    );

    assign s3_shin_valid_i = shin_valid_i;
    assign s3_shin_data_i = shin_data_i[(`SARRAY_LOAD_WIDTH/`SARRAY_H*4)-1:(`SARRAY_LOAD_WIDTH/`SARRAY_H*3)];
    assign sho_valid_o[3] = s3_sho_valid_o;
    assign sho_data_o[(`SARRAY_LOAD_WIDTH/`SARRAY_H*4)-1:(`SARRAY_LOAD_WIDTH/`SARRAY_H*3)] = s3_sho_data_o;



    // -------- shift_reg4

    wire [0:0]                                   s4_shin_valid_i;
    wire [`SARRAY_LOAD_WIDTH/`SARRAY_H-1:0]      s4_shin_data_i;
    wire [0:0]                                   s4_sho_valid_o;
    wire [`SARRAY_LOAD_WIDTH/`SARRAY_H-1:0]      s4_sho_data_o;

    shift_reg #(5) u_shift_reg4 (
        .clk           (clk),
        .rst_n         (rst_n),
        .shin_valid_i  (s4_shin_valid_i),
        .shin_data_i   (s4_shin_data_i),
        .sho_valid_o   (s4_sho_valid_o),
        .sho_data_o    (s4_sho_data_o)
    );

    assign s4_shin_valid_i = shin_valid_i;
    assign s4_shin_data_i = shin_data_i[(`SARRAY_LOAD_WIDTH/`SARRAY_H*5)-1:(`SARRAY_LOAD_WIDTH/`SARRAY_H*4)];
    assign sho_valid_o[4] = s4_sho_valid_o;
    assign sho_data_o[(`SARRAY_LOAD_WIDTH/`SARRAY_H*5)-1:(`SARRAY_LOAD_WIDTH/`SARRAY_H*4)] = s4_sho_data_o;



    // -------- shift_reg5

    wire [0:0]                                   s5_shin_valid_i;
    wire [`SARRAY_LOAD_WIDTH/`SARRAY_H-1:0]      s5_shin_data_i;
    wire [0:0]                                   s5_sho_valid_o;
    wire [`SARRAY_LOAD_WIDTH/`SARRAY_H-1:0]      s5_sho_data_o;

    shift_reg #(6) u_shift_reg5 (
        .clk           (clk),
        .rst_n         (rst_n),
        .shin_valid_i  (s5_shin_valid_i),
        .shin_data_i   (s5_shin_data_i),
        .sho_valid_o   (s5_sho_valid_o),
        .sho_data_o    (s5_sho_data_o)
    );

    assign s5_shin_valid_i = shin_valid_i;
    assign s5_shin_data_i = shin_data_i[(`SARRAY_LOAD_WIDTH/`SARRAY_H*6)-1:(`SARRAY_LOAD_WIDTH/`SARRAY_H*5)];
    assign sho_valid_o[5] = s5_sho_valid_o;
    assign sho_data_o[(`SARRAY_LOAD_WIDTH/`SARRAY_H*6)-1:(`SARRAY_LOAD_WIDTH/`SARRAY_H*5)] = s5_sho_data_o;



    // -------- shift_reg6

    wire [0:0]                                   s6_shin_valid_i;
    wire [`SARRAY_LOAD_WIDTH/`SARRAY_H-1:0]      s6_shin_data_i;
    wire [0:0]                                   s6_sho_valid_o;
    wire [`SARRAY_LOAD_WIDTH/`SARRAY_H-1:0]      s6_sho_data_o;

    shift_reg #(7) u_shift_reg6 (
        .clk           (clk),
        .rst_n         (rst_n),
        .shin_valid_i  (s6_shin_valid_i),
        .shin_data_i   (s6_shin_data_i),
        .sho_valid_o   (s6_sho_valid_o),
        .sho_data_o    (s6_sho_data_o)
    );

    assign s6_shin_valid_i = shin_valid_i;
    assign s6_shin_data_i = shin_data_i[(`SARRAY_LOAD_WIDTH/`SARRAY_H*7)-1:(`SARRAY_LOAD_WIDTH/`SARRAY_H*6)];
    assign sho_valid_o[6] = s6_sho_valid_o;
    assign sho_data_o[(`SARRAY_LOAD_WIDTH/`SARRAY_H*7)-1:(`SARRAY_LOAD_WIDTH/`SARRAY_H*6)] = s6_sho_data_o;



    // -------- shift_reg7

    wire [0:0]                                   s7_shin_valid_i;
    wire [`SARRAY_LOAD_WIDTH/`SARRAY_H-1:0]      s7_shin_data_i;
    wire [0:0]                                   s7_sho_valid_o;
    wire [`SARRAY_LOAD_WIDTH/`SARRAY_H-1:0]      s7_sho_data_o;

    shift_reg #(8) u_shift_reg7 (
        .clk           (clk),
        .rst_n         (rst_n),
        .shin_valid_i  (s7_shin_valid_i),
        .shin_data_i   (s7_shin_data_i),
        .sho_valid_o   (s7_sho_valid_o),
        .sho_data_o    (s7_sho_data_o)
    );

    assign s7_shin_valid_i = shin_valid_i;
    assign s7_shin_data_i = shin_data_i[(`SARRAY_LOAD_WIDTH/`SARRAY_H*8)-1:(`SARRAY_LOAD_WIDTH/`SARRAY_H*7)];
    assign sho_valid_o[7] = s7_sho_valid_o;
    assign sho_data_o[(`SARRAY_LOAD_WIDTH/`SARRAY_H*8)-1:(`SARRAY_LOAD_WIDTH/`SARRAY_H*7)] = s7_sho_data_o;



    // -------- shift_reg8

    wire [0:0]                                   s8_shin_valid_i;
    wire [`SARRAY_LOAD_WIDTH/`SARRAY_H-1:0]      s8_shin_data_i;
    wire [0:0]                                   s8_sho_valid_o;
    wire [`SARRAY_LOAD_WIDTH/`SARRAY_H-1:0]      s8_sho_data_o;

    shift_reg #(9) u_shift_reg8 (
        .clk           (clk),
        .rst_n         (rst_n),
        .shin_valid_i  (s8_shin_valid_i),
        .shin_data_i   (s8_shin_data_i),
        .sho_valid_o   (s8_sho_valid_o),
        .sho_data_o    (s8_sho_data_o)
    );

    assign s8_shin_valid_i = shin_valid_i;
    assign s8_shin_data_i = shin_data_i[(`SARRAY_LOAD_WIDTH/`SARRAY_H*9)-1:(`SARRAY_LOAD_WIDTH/`SARRAY_H*8)];
    assign sho_valid_o[8] = s8_sho_valid_o;
    assign sho_data_o[(`SARRAY_LOAD_WIDTH/`SARRAY_H*9)-1:(`SARRAY_LOAD_WIDTH/`SARRAY_H*8)] = s8_sho_data_o;



    // -------- shift_reg9

    wire [0:0]                                   s9_shin_valid_i;
    wire [`SARRAY_LOAD_WIDTH/`SARRAY_H-1:0]      s9_shin_data_i;
    wire [0:0]                                   s9_sho_valid_o;
    wire [`SARRAY_LOAD_WIDTH/`SARRAY_H-1:0]      s9_sho_data_o;

    shift_reg #(10) u_shift_reg9 (
        .clk           (clk),
        .rst_n         (rst_n),
        .shin_valid_i  (s9_shin_valid_i),
        .shin_data_i   (s9_shin_data_i),
        .sho_valid_o   (s9_sho_valid_o),
        .sho_data_o    (s9_sho_data_o)
    );

    assign s9_shin_valid_i = shin_valid_i;
    assign s9_shin_data_i = shin_data_i[(`SARRAY_LOAD_WIDTH/`SARRAY_H*10)-1:(`SARRAY_LOAD_WIDTH/`SARRAY_H*9)];
    assign sho_valid_o[9] = s9_sho_valid_o;
    assign sho_data_o[(`SARRAY_LOAD_WIDTH/`SARRAY_H*10)-1:(`SARRAY_LOAD_WIDTH/`SARRAY_H*9)] = s9_sho_data_o;



    // -------- shift_reg10

    wire [0:0]                                   s10_shin_valid_i;
    wire [`SARRAY_LOAD_WIDTH/`SARRAY_H-1:0]      s10_shin_data_i;
    wire [0:0]                                   s10_sho_valid_o;
    wire [`SARRAY_LOAD_WIDTH/`SARRAY_H-1:0]      s10_sho_data_o;

    shift_reg #(11) u_shift_reg10 (
        .clk           (clk),
        .rst_n         (rst_n),
        .shin_valid_i  (s10_shin_valid_i),
        .shin_data_i   (s10_shin_data_i),
        .sho_valid_o   (s10_sho_valid_o),
        .sho_data_o    (s10_sho_data_o)
    );

    assign s10_shin_valid_i = shin_valid_i;
    assign s10_shin_data_i = shin_data_i[(`SARRAY_LOAD_WIDTH/`SARRAY_H*11)-1:(`SARRAY_LOAD_WIDTH/`SARRAY_H*10)];
    assign sho_valid_o[10] = s10_sho_valid_o;
    assign sho_data_o[(`SARRAY_LOAD_WIDTH/`SARRAY_H*11)-1:(`SARRAY_LOAD_WIDTH/`SARRAY_H*10)] = s10_sho_data_o;



    // -------- shift_reg11

    wire [0:0]                                   s11_shin_valid_i;
    wire [`SARRAY_LOAD_WIDTH/`SARRAY_H-1:0]      s11_shin_data_i;
    wire [0:0]                                   s11_sho_valid_o;
    wire [`SARRAY_LOAD_WIDTH/`SARRAY_H-1:0]      s11_sho_data_o;

    shift_reg #(12) u_shift_reg11 (
        .clk           (clk),
        .rst_n         (rst_n),
        .shin_valid_i  (s11_shin_valid_i),
        .shin_data_i   (s11_shin_data_i),
        .sho_valid_o   (s11_sho_valid_o),
        .sho_data_o    (s11_sho_data_o)
    );

    assign s11_shin_valid_i = shin_valid_i;
    assign s11_shin_data_i = shin_data_i[(`SARRAY_LOAD_WIDTH/`SARRAY_H*12)-1:(`SARRAY_LOAD_WIDTH/`SARRAY_H*11)];
    assign sho_valid_o[11] = s11_sho_valid_o;
    assign sho_data_o[(`SARRAY_LOAD_WIDTH/`SARRAY_H*12)-1:(`SARRAY_LOAD_WIDTH/`SARRAY_H*11)] = s11_sho_data_o;



    // -------- shift_reg12

    wire [0:0]                                   s12_shin_valid_i;
    wire [`SARRAY_LOAD_WIDTH/`SARRAY_H-1:0]      s12_shin_data_i;
    wire [0:0]                                   s12_sho_valid_o;
    wire [`SARRAY_LOAD_WIDTH/`SARRAY_H-1:0]      s12_sho_data_o;

    shift_reg #(13) u_shift_reg12 (
        .clk           (clk),
        .rst_n         (rst_n),
        .shin_valid_i  (s12_shin_valid_i),
        .shin_data_i   (s12_shin_data_i),
        .sho_valid_o   (s12_sho_valid_o),
        .sho_data_o    (s12_sho_data_o)
    );

    assign s12_shin_valid_i = shin_valid_i;
    assign s12_shin_data_i = shin_data_i[(`SARRAY_LOAD_WIDTH/`SARRAY_H*13)-1:(`SARRAY_LOAD_WIDTH/`SARRAY_H*12)];
    assign sho_valid_o[12] = s12_sho_valid_o;
    assign sho_data_o[(`SARRAY_LOAD_WIDTH/`SARRAY_H*13)-1:(`SARRAY_LOAD_WIDTH/`SARRAY_H*12)] = s12_sho_data_o;



    // -------- shift_reg13

    wire [0:0]                                   s13_shin_valid_i;
    wire [`SARRAY_LOAD_WIDTH/`SARRAY_H-1:0]      s13_shin_data_i;
    wire [0:0]                                   s13_sho_valid_o;
    wire [`SARRAY_LOAD_WIDTH/`SARRAY_H-1:0]      s13_sho_data_o;

    shift_reg #(14) u_shift_reg13 (
        .clk           (clk),
        .rst_n         (rst_n),
        .shin_valid_i  (s13_shin_valid_i),
        .shin_data_i   (s13_shin_data_i),
        .sho_valid_o   (s13_sho_valid_o),
        .sho_data_o    (s13_sho_data_o)
    );

    assign s13_shin_valid_i = shin_valid_i;
    assign s13_shin_data_i = shin_data_i[(`SARRAY_LOAD_WIDTH/`SARRAY_H*14)-1:(`SARRAY_LOAD_WIDTH/`SARRAY_H*13)];
    assign sho_valid_o[13] = s13_sho_valid_o;
    assign sho_data_o[(`SARRAY_LOAD_WIDTH/`SARRAY_H*14)-1:(`SARRAY_LOAD_WIDTH/`SARRAY_H*13)] = s13_sho_data_o;



    // -------- shift_reg14

    wire [0:0]                                   s14_shin_valid_i;
    wire [`SARRAY_LOAD_WIDTH/`SARRAY_H-1:0]      s14_shin_data_i;
    wire [0:0]                                   s14_sho_valid_o;
    wire [`SARRAY_LOAD_WIDTH/`SARRAY_H-1:0]      s14_sho_data_o;

    shift_reg #(15) u_shift_reg14 (
        .clk           (clk),
        .rst_n         (rst_n),
        .shin_valid_i  (s14_shin_valid_i),
        .shin_data_i   (s14_shin_data_i),
        .sho_valid_o   (s14_sho_valid_o),
        .sho_data_o    (s14_sho_data_o)
    );

    assign s14_shin_valid_i = shin_valid_i;
    assign s14_shin_data_i = shin_data_i[(`SARRAY_LOAD_WIDTH/`SARRAY_H*15)-1:(`SARRAY_LOAD_WIDTH/`SARRAY_H*14)];
    assign sho_valid_o[14] = s14_sho_valid_o;
    assign sho_data_o[(`SARRAY_LOAD_WIDTH/`SARRAY_H*15)-1:(`SARRAY_LOAD_WIDTH/`SARRAY_H*14)] = s14_sho_data_o;



    // -------- shift_reg15

    wire [0:0]                                   s15_shin_valid_i;
    wire [`SARRAY_LOAD_WIDTH/`SARRAY_H-1:0]      s15_shin_data_i;
    wire [0:0]                                   s15_sho_valid_o;
    wire [`SARRAY_LOAD_WIDTH/`SARRAY_H-1:0]      s15_sho_data_o;

    shift_reg #(16) u_shift_reg15 (
        .clk           (clk),
        .rst_n         (rst_n),
        .shin_valid_i  (s15_shin_valid_i),
        .shin_data_i   (s15_shin_data_i),
        .sho_valid_o   (s15_sho_valid_o),
        .sho_data_o    (s15_sho_data_o)
    );

    assign s15_shin_valid_i = shin_valid_i;
    assign s15_shin_data_i = shin_data_i[(`SARRAY_LOAD_WIDTH/`SARRAY_H*16)-1:(`SARRAY_LOAD_WIDTH/`SARRAY_H*15)];
    assign sho_valid_o[15] = s15_sho_valid_o;
    assign sho_data_o[(`SARRAY_LOAD_WIDTH/`SARRAY_H*16)-1:(`SARRAY_LOAD_WIDTH/`SARRAY_H*15)] = s15_sho_data_o;



    // -------- shift_reg16

    wire [0:0]                                   s16_shin_valid_i;
    wire [`SARRAY_LOAD_WIDTH/`SARRAY_H-1:0]      s16_shin_data_i;
    wire [0:0]                                   s16_sho_valid_o;
    wire [`SARRAY_LOAD_WIDTH/`SARRAY_H-1:0]      s16_sho_data_o;

    shift_reg #(17) u_shift_reg16 (
        .clk           (clk),
        .rst_n         (rst_n),
        .shin_valid_i  (s16_shin_valid_i),
        .shin_data_i   (s16_shin_data_i),
        .sho_valid_o   (s16_sho_valid_o),
        .sho_data_o    (s16_sho_data_o)
    );

    assign s16_shin_valid_i = shin_valid_i;
    assign s16_shin_data_i = shin_data_i[(`SARRAY_LOAD_WIDTH/`SARRAY_H*17)-1:(`SARRAY_LOAD_WIDTH/`SARRAY_H*16)];
    assign sho_valid_o[16] = s16_sho_valid_o;
    assign sho_data_o[(`SARRAY_LOAD_WIDTH/`SARRAY_H*17)-1:(`SARRAY_LOAD_WIDTH/`SARRAY_H*16)] = s16_sho_data_o;



    // -------- shift_reg17

    wire [0:0]                                   s17_shin_valid_i;
    wire [`SARRAY_LOAD_WIDTH/`SARRAY_H-1:0]      s17_shin_data_i;
    wire [0:0]                                   s17_sho_valid_o;
    wire [`SARRAY_LOAD_WIDTH/`SARRAY_H-1:0]      s17_sho_data_o;

    shift_reg #(18) u_shift_reg17 (
        .clk           (clk),
        .rst_n         (rst_n),
        .shin_valid_i  (s17_shin_valid_i),
        .shin_data_i   (s17_shin_data_i),
        .sho_valid_o   (s17_sho_valid_o),
        .sho_data_o    (s17_sho_data_o)
    );

    assign s17_shin_valid_i = shin_valid_i;
    assign s17_shin_data_i = shin_data_i[(`SARRAY_LOAD_WIDTH/`SARRAY_H*18)-1:(`SARRAY_LOAD_WIDTH/`SARRAY_H*17)];
    assign sho_valid_o[17] = s17_sho_valid_o;
    assign sho_data_o[(`SARRAY_LOAD_WIDTH/`SARRAY_H*18)-1:(`SARRAY_LOAD_WIDTH/`SARRAY_H*17)] = s17_sho_data_o;



    // -------- shift_reg18

    wire [0:0]                                   s18_shin_valid_i;
    wire [`SARRAY_LOAD_WIDTH/`SARRAY_H-1:0]      s18_shin_data_i;
    wire [0:0]                                   s18_sho_valid_o;
    wire [`SARRAY_LOAD_WIDTH/`SARRAY_H-1:0]      s18_sho_data_o;

    shift_reg #(19) u_shift_reg18 (
        .clk           (clk),
        .rst_n         (rst_n),
        .shin_valid_i  (s18_shin_valid_i),
        .shin_data_i   (s18_shin_data_i),
        .sho_valid_o   (s18_sho_valid_o),
        .sho_data_o    (s18_sho_data_o)
    );

    assign s18_shin_valid_i = shin_valid_i;
    assign s18_shin_data_i = shin_data_i[(`SARRAY_LOAD_WIDTH/`SARRAY_H*19)-1:(`SARRAY_LOAD_WIDTH/`SARRAY_H*18)];
    assign sho_valid_o[18] = s18_sho_valid_o;
    assign sho_data_o[(`SARRAY_LOAD_WIDTH/`SARRAY_H*19)-1:(`SARRAY_LOAD_WIDTH/`SARRAY_H*18)] = s18_sho_data_o;



    // -------- shift_reg19

    wire [0:0]                                   s19_shin_valid_i;
    wire [`SARRAY_LOAD_WIDTH/`SARRAY_H-1:0]      s19_shin_data_i;
    wire [0:0]                                   s19_sho_valid_o;
    wire [`SARRAY_LOAD_WIDTH/`SARRAY_H-1:0]      s19_sho_data_o;

    shift_reg #(20) u_shift_reg19 (
        .clk           (clk),
        .rst_n         (rst_n),
        .shin_valid_i  (s19_shin_valid_i),
        .shin_data_i   (s19_shin_data_i),
        .sho_valid_o   (s19_sho_valid_o),
        .sho_data_o    (s19_sho_data_o)
    );

    assign s19_shin_valid_i = shin_valid_i;
    assign s19_shin_data_i = shin_data_i[(`SARRAY_LOAD_WIDTH/`SARRAY_H*20)-1:(`SARRAY_LOAD_WIDTH/`SARRAY_H*19)];
    assign sho_valid_o[19] = s19_sho_valid_o;
    assign sho_data_o[(`SARRAY_LOAD_WIDTH/`SARRAY_H*20)-1:(`SARRAY_LOAD_WIDTH/`SARRAY_H*19)] = s19_sho_data_o;



    // -------- shift_reg20

    wire [0:0]                                   s20_shin_valid_i;
    wire [`SARRAY_LOAD_WIDTH/`SARRAY_H-1:0]      s20_shin_data_i;
    wire [0:0]                                   s20_sho_valid_o;
    wire [`SARRAY_LOAD_WIDTH/`SARRAY_H-1:0]      s20_sho_data_o;

    shift_reg #(21) u_shift_reg20 (
        .clk           (clk),
        .rst_n         (rst_n),
        .shin_valid_i  (s20_shin_valid_i),
        .shin_data_i   (s20_shin_data_i),
        .sho_valid_o   (s20_sho_valid_o),
        .sho_data_o    (s20_sho_data_o)
    );

    assign s20_shin_valid_i = shin_valid_i;
    assign s20_shin_data_i = shin_data_i[(`SARRAY_LOAD_WIDTH/`SARRAY_H*21)-1:(`SARRAY_LOAD_WIDTH/`SARRAY_H*20)];
    assign sho_valid_o[20] = s20_sho_valid_o;
    assign sho_data_o[(`SARRAY_LOAD_WIDTH/`SARRAY_H*21)-1:(`SARRAY_LOAD_WIDTH/`SARRAY_H*20)] = s20_sho_data_o;



    // -------- shift_reg21

    wire [0:0]                                   s21_shin_valid_i;
    wire [`SARRAY_LOAD_WIDTH/`SARRAY_H-1:0]      s21_shin_data_i;
    wire [0:0]                                   s21_sho_valid_o;
    wire [`SARRAY_LOAD_WIDTH/`SARRAY_H-1:0]      s21_sho_data_o;

    shift_reg #(22) u_shift_reg21 (
        .clk           (clk),
        .rst_n         (rst_n),
        .shin_valid_i  (s21_shin_valid_i),
        .shin_data_i   (s21_shin_data_i),
        .sho_valid_o   (s21_sho_valid_o),
        .sho_data_o    (s21_sho_data_o)
    );

    assign s21_shin_valid_i = shin_valid_i;
    assign s21_shin_data_i = shin_data_i[(`SARRAY_LOAD_WIDTH/`SARRAY_H*22)-1:(`SARRAY_LOAD_WIDTH/`SARRAY_H*21)];
    assign sho_valid_o[21] = s21_sho_valid_o;
    assign sho_data_o[(`SARRAY_LOAD_WIDTH/`SARRAY_H*22)-1:(`SARRAY_LOAD_WIDTH/`SARRAY_H*21)] = s21_sho_data_o;



    // -------- shift_reg22

    wire [0:0]                                   s22_shin_valid_i;
    wire [`SARRAY_LOAD_WIDTH/`SARRAY_H-1:0]      s22_shin_data_i;
    wire [0:0]                                   s22_sho_valid_o;
    wire [`SARRAY_LOAD_WIDTH/`SARRAY_H-1:0]      s22_sho_data_o;

    shift_reg #(23) u_shift_reg22 (
        .clk           (clk),
        .rst_n         (rst_n),
        .shin_valid_i  (s22_shin_valid_i),
        .shin_data_i   (s22_shin_data_i),
        .sho_valid_o   (s22_sho_valid_o),
        .sho_data_o    (s22_sho_data_o)
    );

    assign s22_shin_valid_i = shin_valid_i;
    assign s22_shin_data_i = shin_data_i[(`SARRAY_LOAD_WIDTH/`SARRAY_H*23)-1:(`SARRAY_LOAD_WIDTH/`SARRAY_H*22)];
    assign sho_valid_o[22] = s22_sho_valid_o;
    assign sho_data_o[(`SARRAY_LOAD_WIDTH/`SARRAY_H*23)-1:(`SARRAY_LOAD_WIDTH/`SARRAY_H*22)] = s22_sho_data_o;



    // -------- shift_reg23

    wire [0:0]                                   s23_shin_valid_i;
    wire [`SARRAY_LOAD_WIDTH/`SARRAY_H-1:0]      s23_shin_data_i;
    wire [0:0]                                   s23_sho_valid_o;
    wire [`SARRAY_LOAD_WIDTH/`SARRAY_H-1:0]      s23_sho_data_o;

    shift_reg #(24) u_shift_reg23 (
        .clk           (clk),
        .rst_n         (rst_n),
        .shin_valid_i  (s23_shin_valid_i),
        .shin_data_i   (s23_shin_data_i),
        .sho_valid_o   (s23_sho_valid_o),
        .sho_data_o    (s23_sho_data_o)
    );

    assign s23_shin_valid_i = shin_valid_i;
    assign s23_shin_data_i = shin_data_i[(`SARRAY_LOAD_WIDTH/`SARRAY_H*24)-1:(`SARRAY_LOAD_WIDTH/`SARRAY_H*23)];
    assign sho_valid_o[23] = s23_sho_valid_o;
    assign sho_data_o[(`SARRAY_LOAD_WIDTH/`SARRAY_H*24)-1:(`SARRAY_LOAD_WIDTH/`SARRAY_H*23)] = s23_sho_data_o;



    // -------- shift_reg24

    wire [0:0]                                   s24_shin_valid_i;
    wire [`SARRAY_LOAD_WIDTH/`SARRAY_H-1:0]      s24_shin_data_i;
    wire [0:0]                                   s24_sho_valid_o;
    wire [`SARRAY_LOAD_WIDTH/`SARRAY_H-1:0]      s24_sho_data_o;

    shift_reg #(25) u_shift_reg24 (
        .clk           (clk),
        .rst_n         (rst_n),
        .shin_valid_i  (s24_shin_valid_i),
        .shin_data_i   (s24_shin_data_i),
        .sho_valid_o   (s24_sho_valid_o),
        .sho_data_o    (s24_sho_data_o)
    );

    assign s24_shin_valid_i = shin_valid_i;
    assign s24_shin_data_i = shin_data_i[(`SARRAY_LOAD_WIDTH/`SARRAY_H*25)-1:(`SARRAY_LOAD_WIDTH/`SARRAY_H*24)];
    assign sho_valid_o[24] = s24_sho_valid_o;
    assign sho_data_o[(`SARRAY_LOAD_WIDTH/`SARRAY_H*25)-1:(`SARRAY_LOAD_WIDTH/`SARRAY_H*24)] = s24_sho_data_o;



    // -------- shift_reg25

    wire [0:0]                                   s25_shin_valid_i;
    wire [`SARRAY_LOAD_WIDTH/`SARRAY_H-1:0]      s25_shin_data_i;
    wire [0:0]                                   s25_sho_valid_o;
    wire [`SARRAY_LOAD_WIDTH/`SARRAY_H-1:0]      s25_sho_data_o;

    shift_reg #(26) u_shift_reg25 (
        .clk           (clk),
        .rst_n         (rst_n),
        .shin_valid_i  (s25_shin_valid_i),
        .shin_data_i   (s25_shin_data_i),
        .sho_valid_o   (s25_sho_valid_o),
        .sho_data_o    (s25_sho_data_o)
    );

    assign s25_shin_valid_i = shin_valid_i;
    assign s25_shin_data_i = shin_data_i[(`SARRAY_LOAD_WIDTH/`SARRAY_H*26)-1:(`SARRAY_LOAD_WIDTH/`SARRAY_H*25)];
    assign sho_valid_o[25] = s25_sho_valid_o;
    assign sho_data_o[(`SARRAY_LOAD_WIDTH/`SARRAY_H*26)-1:(`SARRAY_LOAD_WIDTH/`SARRAY_H*25)] = s25_sho_data_o;



    // -------- shift_reg26

    wire [0:0]                                   s26_shin_valid_i;
    wire [`SARRAY_LOAD_WIDTH/`SARRAY_H-1:0]      s26_shin_data_i;
    wire [0:0]                                   s26_sho_valid_o;
    wire [`SARRAY_LOAD_WIDTH/`SARRAY_H-1:0]      s26_sho_data_o;

    shift_reg #(27) u_shift_reg26 (
        .clk           (clk),
        .rst_n         (rst_n),
        .shin_valid_i  (s26_shin_valid_i),
        .shin_data_i   (s26_shin_data_i),
        .sho_valid_o   (s26_sho_valid_o),
        .sho_data_o    (s26_sho_data_o)
    );

    assign s26_shin_valid_i = shin_valid_i;
    assign s26_shin_data_i = shin_data_i[(`SARRAY_LOAD_WIDTH/`SARRAY_H*27)-1:(`SARRAY_LOAD_WIDTH/`SARRAY_H*26)];
    assign sho_valid_o[26] = s26_sho_valid_o;
    assign sho_data_o[(`SARRAY_LOAD_WIDTH/`SARRAY_H*27)-1:(`SARRAY_LOAD_WIDTH/`SARRAY_H*26)] = s26_sho_data_o;



    // -------- shift_reg27

    wire [0:0]                                   s27_shin_valid_i;
    wire [`SARRAY_LOAD_WIDTH/`SARRAY_H-1:0]      s27_shin_data_i;
    wire [0:0]                                   s27_sho_valid_o;
    wire [`SARRAY_LOAD_WIDTH/`SARRAY_H-1:0]      s27_sho_data_o;

    shift_reg #(28) u_shift_reg27 (
        .clk           (clk),
        .rst_n         (rst_n),
        .shin_valid_i  (s27_shin_valid_i),
        .shin_data_i   (s27_shin_data_i),
        .sho_valid_o   (s27_sho_valid_o),
        .sho_data_o    (s27_sho_data_o)
    );

    assign s27_shin_valid_i = shin_valid_i;
    assign s27_shin_data_i = shin_data_i[(`SARRAY_LOAD_WIDTH/`SARRAY_H*28)-1:(`SARRAY_LOAD_WIDTH/`SARRAY_H*27)];
    assign sho_valid_o[27] = s27_sho_valid_o;
    assign sho_data_o[(`SARRAY_LOAD_WIDTH/`SARRAY_H*28)-1:(`SARRAY_LOAD_WIDTH/`SARRAY_H*27)] = s27_sho_data_o;



    // -------- shift_reg28

    wire [0:0]                                   s28_shin_valid_i;
    wire [`SARRAY_LOAD_WIDTH/`SARRAY_H-1:0]      s28_shin_data_i;
    wire [0:0]                                   s28_sho_valid_o;
    wire [`SARRAY_LOAD_WIDTH/`SARRAY_H-1:0]      s28_sho_data_o;

    shift_reg #(29) u_shift_reg28 (
        .clk           (clk),
        .rst_n         (rst_n),
        .shin_valid_i  (s28_shin_valid_i),
        .shin_data_i   (s28_shin_data_i),
        .sho_valid_o   (s28_sho_valid_o),
        .sho_data_o    (s28_sho_data_o)
    );

    assign s28_shin_valid_i = shin_valid_i;
    assign s28_shin_data_i = shin_data_i[(`SARRAY_LOAD_WIDTH/`SARRAY_H*29)-1:(`SARRAY_LOAD_WIDTH/`SARRAY_H*28)];
    assign sho_valid_o[28] = s28_sho_valid_o;
    assign sho_data_o[(`SARRAY_LOAD_WIDTH/`SARRAY_H*29)-1:(`SARRAY_LOAD_WIDTH/`SARRAY_H*28)] = s28_sho_data_o;



    // -------- shift_reg29

    wire [0:0]                                   s29_shin_valid_i;
    wire [`SARRAY_LOAD_WIDTH/`SARRAY_H-1:0]      s29_shin_data_i;
    wire [0:0]                                   s29_sho_valid_o;
    wire [`SARRAY_LOAD_WIDTH/`SARRAY_H-1:0]      s29_sho_data_o;

    shift_reg #(30) u_shift_reg29 (
        .clk           (clk),
        .rst_n         (rst_n),
        .shin_valid_i  (s29_shin_valid_i),
        .shin_data_i   (s29_shin_data_i),
        .sho_valid_o   (s29_sho_valid_o),
        .sho_data_o    (s29_sho_data_o)
    );

    assign s29_shin_valid_i = shin_valid_i;
    assign s29_shin_data_i = shin_data_i[(`SARRAY_LOAD_WIDTH/`SARRAY_H*30)-1:(`SARRAY_LOAD_WIDTH/`SARRAY_H*29)];
    assign sho_valid_o[29] = s29_sho_valid_o;
    assign sho_data_o[(`SARRAY_LOAD_WIDTH/`SARRAY_H*30)-1:(`SARRAY_LOAD_WIDTH/`SARRAY_H*29)] = s29_sho_data_o;



    // -------- shift_reg30

    wire [0:0]                                   s30_shin_valid_i;
    wire [`SARRAY_LOAD_WIDTH/`SARRAY_H-1:0]      s30_shin_data_i;
    wire [0:0]                                   s30_sho_valid_o;
    wire [`SARRAY_LOAD_WIDTH/`SARRAY_H-1:0]      s30_sho_data_o;

    shift_reg #(31) u_shift_reg30 (
        .clk           (clk),
        .rst_n         (rst_n),
        .shin_valid_i  (s30_shin_valid_i),
        .shin_data_i   (s30_shin_data_i),
        .sho_valid_o   (s30_sho_valid_o),
        .sho_data_o    (s30_sho_data_o)
    );

    assign s30_shin_valid_i = shin_valid_i;
    assign s30_shin_data_i = shin_data_i[(`SARRAY_LOAD_WIDTH/`SARRAY_H*31)-1:(`SARRAY_LOAD_WIDTH/`SARRAY_H*30)];
    assign sho_valid_o[30] = s30_sho_valid_o;
    assign sho_data_o[(`SARRAY_LOAD_WIDTH/`SARRAY_H*31)-1:(`SARRAY_LOAD_WIDTH/`SARRAY_H*30)] = s30_sho_data_o;



    // -------- shift_reg31

    wire [0:0]                                   s31_shin_valid_i;
    wire [`SARRAY_LOAD_WIDTH/`SARRAY_H-1:0]      s31_shin_data_i;
    wire [0:0]                                   s31_sho_valid_o;
    wire [`SARRAY_LOAD_WIDTH/`SARRAY_H-1:0]      s31_sho_data_o;

    shift_reg #(32) u_shift_reg31 (
        .clk           (clk),
        .rst_n         (rst_n),
        .shin_valid_i  (s31_shin_valid_i),
        .shin_data_i   (s31_shin_data_i),
        .sho_valid_o   (s31_sho_valid_o),
        .sho_data_o    (s31_sho_data_o)
    );

    assign s31_shin_valid_i = shin_valid_i;
    assign s31_shin_data_i = shin_data_i[(`SARRAY_LOAD_WIDTH/`SARRAY_H*32)-1:(`SARRAY_LOAD_WIDTH/`SARRAY_H*31)];
    assign sho_valid_o[31] = s31_sho_valid_o;
    assign sho_data_o[(`SARRAY_LOAD_WIDTH/`SARRAY_H*32)-1:(`SARRAY_LOAD_WIDTH/`SARRAY_H*31)] = s31_sho_data_o;



    // -------- shift_reg32

    wire [0:0]                                   s32_shin_valid_i;
    wire [`SARRAY_LOAD_WIDTH/`SARRAY_H-1:0]      s32_shin_data_i;
    wire [0:0]                                   s32_sho_valid_o;
    wire [`SARRAY_LOAD_WIDTH/`SARRAY_H-1:0]      s32_sho_data_o;

    shift_reg #(33) u_shift_reg32 (
        .clk           (clk),
        .rst_n         (rst_n),
        .shin_valid_i  (s32_shin_valid_i),
        .shin_data_i   (s32_shin_data_i),
        .sho_valid_o   (s32_sho_valid_o),
        .sho_data_o    (s32_sho_data_o)
    );

    assign s32_shin_valid_i = shin_valid_i;
    assign s32_shin_data_i = shin_data_i[(`SARRAY_LOAD_WIDTH/`SARRAY_H*33)-1:(`SARRAY_LOAD_WIDTH/`SARRAY_H*32)];
    assign sho_valid_o[32] = s32_sho_valid_o;
    assign sho_data_o[(`SARRAY_LOAD_WIDTH/`SARRAY_H*33)-1:(`SARRAY_LOAD_WIDTH/`SARRAY_H*32)] = s32_sho_data_o;



    // -------- shift_reg33

    wire [0:0]                                   s33_shin_valid_i;
    wire [`SARRAY_LOAD_WIDTH/`SARRAY_H-1:0]      s33_shin_data_i;
    wire [0:0]                                   s33_sho_valid_o;
    wire [`SARRAY_LOAD_WIDTH/`SARRAY_H-1:0]      s33_sho_data_o;

    shift_reg #(34) u_shift_reg33 (
        .clk           (clk),
        .rst_n         (rst_n),
        .shin_valid_i  (s33_shin_valid_i),
        .shin_data_i   (s33_shin_data_i),
        .sho_valid_o   (s33_sho_valid_o),
        .sho_data_o    (s33_sho_data_o)
    );

    assign s33_shin_valid_i = shin_valid_i;
    assign s33_shin_data_i = shin_data_i[(`SARRAY_LOAD_WIDTH/`SARRAY_H*34)-1:(`SARRAY_LOAD_WIDTH/`SARRAY_H*33)];
    assign sho_valid_o[33] = s33_sho_valid_o;
    assign sho_data_o[(`SARRAY_LOAD_WIDTH/`SARRAY_H*34)-1:(`SARRAY_LOAD_WIDTH/`SARRAY_H*33)] = s33_sho_data_o;



    // -------- shift_reg34

    wire [0:0]                                   s34_shin_valid_i;
    wire [`SARRAY_LOAD_WIDTH/`SARRAY_H-1:0]      s34_shin_data_i;
    wire [0:0]                                   s34_sho_valid_o;
    wire [`SARRAY_LOAD_WIDTH/`SARRAY_H-1:0]      s34_sho_data_o;

    shift_reg #(35) u_shift_reg34 (
        .clk           (clk),
        .rst_n         (rst_n),
        .shin_valid_i  (s34_shin_valid_i),
        .shin_data_i   (s34_shin_data_i),
        .sho_valid_o   (s34_sho_valid_o),
        .sho_data_o    (s34_sho_data_o)
    );

    assign s34_shin_valid_i = shin_valid_i;
    assign s34_shin_data_i = shin_data_i[(`SARRAY_LOAD_WIDTH/`SARRAY_H*35)-1:(`SARRAY_LOAD_WIDTH/`SARRAY_H*34)];
    assign sho_valid_o[34] = s34_sho_valid_o;
    assign sho_data_o[(`SARRAY_LOAD_WIDTH/`SARRAY_H*35)-1:(`SARRAY_LOAD_WIDTH/`SARRAY_H*34)] = s34_sho_data_o;



    // -------- shift_reg35

    wire [0:0]                                   s35_shin_valid_i;
    wire [`SARRAY_LOAD_WIDTH/`SARRAY_H-1:0]      s35_shin_data_i;
    wire [0:0]                                   s35_sho_valid_o;
    wire [`SARRAY_LOAD_WIDTH/`SARRAY_H-1:0]      s35_sho_data_o;

    shift_reg #(36) u_shift_reg35 (
        .clk           (clk),
        .rst_n         (rst_n),
        .shin_valid_i  (s35_shin_valid_i),
        .shin_data_i   (s35_shin_data_i),
        .sho_valid_o   (s35_sho_valid_o),
        .sho_data_o    (s35_sho_data_o)
    );

    assign s35_shin_valid_i = shin_valid_i;
    assign s35_shin_data_i = shin_data_i[(`SARRAY_LOAD_WIDTH/`SARRAY_H*36)-1:(`SARRAY_LOAD_WIDTH/`SARRAY_H*35)];
    assign sho_valid_o[35] = s35_sho_valid_o;
    assign sho_data_o[(`SARRAY_LOAD_WIDTH/`SARRAY_H*36)-1:(`SARRAY_LOAD_WIDTH/`SARRAY_H*35)] = s35_sho_data_o;



    // -------- shift_reg36

    wire [0:0]                                   s36_shin_valid_i;
    wire [`SARRAY_LOAD_WIDTH/`SARRAY_H-1:0]      s36_shin_data_i;
    wire [0:0]                                   s36_sho_valid_o;
    wire [`SARRAY_LOAD_WIDTH/`SARRAY_H-1:0]      s36_sho_data_o;

    shift_reg #(37) u_shift_reg36 (
        .clk           (clk),
        .rst_n         (rst_n),
        .shin_valid_i  (s36_shin_valid_i),
        .shin_data_i   (s36_shin_data_i),
        .sho_valid_o   (s36_sho_valid_o),
        .sho_data_o    (s36_sho_data_o)
    );

    assign s36_shin_valid_i = shin_valid_i;
    assign s36_shin_data_i = shin_data_i[(`SARRAY_LOAD_WIDTH/`SARRAY_H*37)-1:(`SARRAY_LOAD_WIDTH/`SARRAY_H*36)];
    assign sho_valid_o[36] = s36_sho_valid_o;
    assign sho_data_o[(`SARRAY_LOAD_WIDTH/`SARRAY_H*37)-1:(`SARRAY_LOAD_WIDTH/`SARRAY_H*36)] = s36_sho_data_o;



    // -------- shift_reg37

    wire [0:0]                                   s37_shin_valid_i;
    wire [`SARRAY_LOAD_WIDTH/`SARRAY_H-1:0]      s37_shin_data_i;
    wire [0:0]                                   s37_sho_valid_o;
    wire [`SARRAY_LOAD_WIDTH/`SARRAY_H-1:0]      s37_sho_data_o;

    shift_reg #(38) u_shift_reg37 (
        .clk           (clk),
        .rst_n         (rst_n),
        .shin_valid_i  (s37_shin_valid_i),
        .shin_data_i   (s37_shin_data_i),
        .sho_valid_o   (s37_sho_valid_o),
        .sho_data_o    (s37_sho_data_o)
    );

    assign s37_shin_valid_i = shin_valid_i;
    assign s37_shin_data_i = shin_data_i[(`SARRAY_LOAD_WIDTH/`SARRAY_H*38)-1:(`SARRAY_LOAD_WIDTH/`SARRAY_H*37)];
    assign sho_valid_o[37] = s37_sho_valid_o;
    assign sho_data_o[(`SARRAY_LOAD_WIDTH/`SARRAY_H*38)-1:(`SARRAY_LOAD_WIDTH/`SARRAY_H*37)] = s37_sho_data_o;



    // -------- shift_reg38

    wire [0:0]                                   s38_shin_valid_i;
    wire [`SARRAY_LOAD_WIDTH/`SARRAY_H-1:0]      s38_shin_data_i;
    wire [0:0]                                   s38_sho_valid_o;
    wire [`SARRAY_LOAD_WIDTH/`SARRAY_H-1:0]      s38_sho_data_o;

    shift_reg #(39) u_shift_reg38 (
        .clk           (clk),
        .rst_n         (rst_n),
        .shin_valid_i  (s38_shin_valid_i),
        .shin_data_i   (s38_shin_data_i),
        .sho_valid_o   (s38_sho_valid_o),
        .sho_data_o    (s38_sho_data_o)
    );

    assign s38_shin_valid_i = shin_valid_i;
    assign s38_shin_data_i = shin_data_i[(`SARRAY_LOAD_WIDTH/`SARRAY_H*39)-1:(`SARRAY_LOAD_WIDTH/`SARRAY_H*38)];
    assign sho_valid_o[38] = s38_sho_valid_o;
    assign sho_data_o[(`SARRAY_LOAD_WIDTH/`SARRAY_H*39)-1:(`SARRAY_LOAD_WIDTH/`SARRAY_H*38)] = s38_sho_data_o;



    // -------- shift_reg39

    wire [0:0]                                   s39_shin_valid_i;
    wire [`SARRAY_LOAD_WIDTH/`SARRAY_H-1:0]      s39_shin_data_i;
    wire [0:0]                                   s39_sho_valid_o;
    wire [`SARRAY_LOAD_WIDTH/`SARRAY_H-1:0]      s39_sho_data_o;

    shift_reg #(40) u_shift_reg39 (
        .clk           (clk),
        .rst_n         (rst_n),
        .shin_valid_i  (s39_shin_valid_i),
        .shin_data_i   (s39_shin_data_i),
        .sho_valid_o   (s39_sho_valid_o),
        .sho_data_o    (s39_sho_data_o)
    );

    assign s39_shin_valid_i = shin_valid_i;
    assign s39_shin_data_i = shin_data_i[(`SARRAY_LOAD_WIDTH/`SARRAY_H*40)-1:(`SARRAY_LOAD_WIDTH/`SARRAY_H*39)];
    assign sho_valid_o[39] = s39_sho_valid_o;
    assign sho_data_o[(`SARRAY_LOAD_WIDTH/`SARRAY_H*40)-1:(`SARRAY_LOAD_WIDTH/`SARRAY_H*39)] = s39_sho_data_o;



    // -------- shift_reg40

    wire [0:0]                                   s40_shin_valid_i;
    wire [`SARRAY_LOAD_WIDTH/`SARRAY_H-1:0]      s40_shin_data_i;
    wire [0:0]                                   s40_sho_valid_o;
    wire [`SARRAY_LOAD_WIDTH/`SARRAY_H-1:0]      s40_sho_data_o;

    shift_reg #(41) u_shift_reg40 (
        .clk           (clk),
        .rst_n         (rst_n),
        .shin_valid_i  (s40_shin_valid_i),
        .shin_data_i   (s40_shin_data_i),
        .sho_valid_o   (s40_sho_valid_o),
        .sho_data_o    (s40_sho_data_o)
    );

    assign s40_shin_valid_i = shin_valid_i;
    assign s40_shin_data_i = shin_data_i[(`SARRAY_LOAD_WIDTH/`SARRAY_H*41)-1:(`SARRAY_LOAD_WIDTH/`SARRAY_H*40)];
    assign sho_valid_o[40] = s40_sho_valid_o;
    assign sho_data_o[(`SARRAY_LOAD_WIDTH/`SARRAY_H*41)-1:(`SARRAY_LOAD_WIDTH/`SARRAY_H*40)] = s40_sho_data_o;



    // -------- shift_reg41

    wire [0:0]                                   s41_shin_valid_i;
    wire [`SARRAY_LOAD_WIDTH/`SARRAY_H-1:0]      s41_shin_data_i;
    wire [0:0]                                   s41_sho_valid_o;
    wire [`SARRAY_LOAD_WIDTH/`SARRAY_H-1:0]      s41_sho_data_o;

    shift_reg #(42) u_shift_reg41 (
        .clk           (clk),
        .rst_n         (rst_n),
        .shin_valid_i  (s41_shin_valid_i),
        .shin_data_i   (s41_shin_data_i),
        .sho_valid_o   (s41_sho_valid_o),
        .sho_data_o    (s41_sho_data_o)
    );

    assign s41_shin_valid_i = shin_valid_i;
    assign s41_shin_data_i = shin_data_i[(`SARRAY_LOAD_WIDTH/`SARRAY_H*42)-1:(`SARRAY_LOAD_WIDTH/`SARRAY_H*41)];
    assign sho_valid_o[41] = s41_sho_valid_o;
    assign sho_data_o[(`SARRAY_LOAD_WIDTH/`SARRAY_H*42)-1:(`SARRAY_LOAD_WIDTH/`SARRAY_H*41)] = s41_sho_data_o;



    // -------- shift_reg42

    wire [0:0]                                   s42_shin_valid_i;
    wire [`SARRAY_LOAD_WIDTH/`SARRAY_H-1:0]      s42_shin_data_i;
    wire [0:0]                                   s42_sho_valid_o;
    wire [`SARRAY_LOAD_WIDTH/`SARRAY_H-1:0]      s42_sho_data_o;

    shift_reg #(43) u_shift_reg42 (
        .clk           (clk),
        .rst_n         (rst_n),
        .shin_valid_i  (s42_shin_valid_i),
        .shin_data_i   (s42_shin_data_i),
        .sho_valid_o   (s42_sho_valid_o),
        .sho_data_o    (s42_sho_data_o)
    );

    assign s42_shin_valid_i = shin_valid_i;
    assign s42_shin_data_i = shin_data_i[(`SARRAY_LOAD_WIDTH/`SARRAY_H*43)-1:(`SARRAY_LOAD_WIDTH/`SARRAY_H*42)];
    assign sho_valid_o[42] = s42_sho_valid_o;
    assign sho_data_o[(`SARRAY_LOAD_WIDTH/`SARRAY_H*43)-1:(`SARRAY_LOAD_WIDTH/`SARRAY_H*42)] = s42_sho_data_o;



    // -------- shift_reg43

    wire [0:0]                                   s43_shin_valid_i;
    wire [`SARRAY_LOAD_WIDTH/`SARRAY_H-1:0]      s43_shin_data_i;
    wire [0:0]                                   s43_sho_valid_o;
    wire [`SARRAY_LOAD_WIDTH/`SARRAY_H-1:0]      s43_sho_data_o;

    shift_reg #(44) u_shift_reg43 (
        .clk           (clk),
        .rst_n         (rst_n),
        .shin_valid_i  (s43_shin_valid_i),
        .shin_data_i   (s43_shin_data_i),
        .sho_valid_o   (s43_sho_valid_o),
        .sho_data_o    (s43_sho_data_o)
    );

    assign s43_shin_valid_i = shin_valid_i;
    assign s43_shin_data_i = shin_data_i[(`SARRAY_LOAD_WIDTH/`SARRAY_H*44)-1:(`SARRAY_LOAD_WIDTH/`SARRAY_H*43)];
    assign sho_valid_o[43] = s43_sho_valid_o;
    assign sho_data_o[(`SARRAY_LOAD_WIDTH/`SARRAY_H*44)-1:(`SARRAY_LOAD_WIDTH/`SARRAY_H*43)] = s43_sho_data_o;



    // -------- shift_reg44

    wire [0:0]                                   s44_shin_valid_i;
    wire [`SARRAY_LOAD_WIDTH/`SARRAY_H-1:0]      s44_shin_data_i;
    wire [0:0]                                   s44_sho_valid_o;
    wire [`SARRAY_LOAD_WIDTH/`SARRAY_H-1:0]      s44_sho_data_o;

    shift_reg #(45) u_shift_reg44 (
        .clk           (clk),
        .rst_n         (rst_n),
        .shin_valid_i  (s44_shin_valid_i),
        .shin_data_i   (s44_shin_data_i),
        .sho_valid_o   (s44_sho_valid_o),
        .sho_data_o    (s44_sho_data_o)
    );

    assign s44_shin_valid_i = shin_valid_i;
    assign s44_shin_data_i = shin_data_i[(`SARRAY_LOAD_WIDTH/`SARRAY_H*45)-1:(`SARRAY_LOAD_WIDTH/`SARRAY_H*44)];
    assign sho_valid_o[44] = s44_sho_valid_o;
    assign sho_data_o[(`SARRAY_LOAD_WIDTH/`SARRAY_H*45)-1:(`SARRAY_LOAD_WIDTH/`SARRAY_H*44)] = s44_sho_data_o;



    // -------- shift_reg45

    wire [0:0]                                   s45_shin_valid_i;
    wire [`SARRAY_LOAD_WIDTH/`SARRAY_H-1:0]      s45_shin_data_i;
    wire [0:0]                                   s45_sho_valid_o;
    wire [`SARRAY_LOAD_WIDTH/`SARRAY_H-1:0]      s45_sho_data_o;

    shift_reg #(46) u_shift_reg45 (
        .clk           (clk),
        .rst_n         (rst_n),
        .shin_valid_i  (s45_shin_valid_i),
        .shin_data_i   (s45_shin_data_i),
        .sho_valid_o   (s45_sho_valid_o),
        .sho_data_o    (s45_sho_data_o)
    );

    assign s45_shin_valid_i = shin_valid_i;
    assign s45_shin_data_i = shin_data_i[(`SARRAY_LOAD_WIDTH/`SARRAY_H*46)-1:(`SARRAY_LOAD_WIDTH/`SARRAY_H*45)];
    assign sho_valid_o[45] = s45_sho_valid_o;
    assign sho_data_o[(`SARRAY_LOAD_WIDTH/`SARRAY_H*46)-1:(`SARRAY_LOAD_WIDTH/`SARRAY_H*45)] = s45_sho_data_o;



    // -------- shift_reg46

    wire [0:0]                                   s46_shin_valid_i;
    wire [`SARRAY_LOAD_WIDTH/`SARRAY_H-1:0]      s46_shin_data_i;
    wire [0:0]                                   s46_sho_valid_o;
    wire [`SARRAY_LOAD_WIDTH/`SARRAY_H-1:0]      s46_sho_data_o;

    shift_reg #(47) u_shift_reg46 (
        .clk           (clk),
        .rst_n         (rst_n),
        .shin_valid_i  (s46_shin_valid_i),
        .shin_data_i   (s46_shin_data_i),
        .sho_valid_o   (s46_sho_valid_o),
        .sho_data_o    (s46_sho_data_o)
    );

    assign s46_shin_valid_i = shin_valid_i;
    assign s46_shin_data_i = shin_data_i[(`SARRAY_LOAD_WIDTH/`SARRAY_H*47)-1:(`SARRAY_LOAD_WIDTH/`SARRAY_H*46)];
    assign sho_valid_o[46] = s46_sho_valid_o;
    assign sho_data_o[(`SARRAY_LOAD_WIDTH/`SARRAY_H*47)-1:(`SARRAY_LOAD_WIDTH/`SARRAY_H*46)] = s46_sho_data_o;



    // -------- shift_reg47

    wire [0:0]                                   s47_shin_valid_i;
    wire [`SARRAY_LOAD_WIDTH/`SARRAY_H-1:0]      s47_shin_data_i;
    wire [0:0]                                   s47_sho_valid_o;
    wire [`SARRAY_LOAD_WIDTH/`SARRAY_H-1:0]      s47_sho_data_o;

    shift_reg #(48) u_shift_reg47 (
        .clk           (clk),
        .rst_n         (rst_n),
        .shin_valid_i  (s47_shin_valid_i),
        .shin_data_i   (s47_shin_data_i),
        .sho_valid_o   (s47_sho_valid_o),
        .sho_data_o    (s47_sho_data_o)
    );

    assign s47_shin_valid_i = shin_valid_i;
    assign s47_shin_data_i = shin_data_i[(`SARRAY_LOAD_WIDTH/`SARRAY_H*48)-1:(`SARRAY_LOAD_WIDTH/`SARRAY_H*47)];
    assign sho_valid_o[47] = s47_sho_valid_o;
    assign sho_data_o[(`SARRAY_LOAD_WIDTH/`SARRAY_H*48)-1:(`SARRAY_LOAD_WIDTH/`SARRAY_H*47)] = s47_sho_data_o;



    // -------- shift_reg48

    wire [0:0]                                   s48_shin_valid_i;
    wire [`SARRAY_LOAD_WIDTH/`SARRAY_H-1:0]      s48_shin_data_i;
    wire [0:0]                                   s48_sho_valid_o;
    wire [`SARRAY_LOAD_WIDTH/`SARRAY_H-1:0]      s48_sho_data_o;

    shift_reg #(49) u_shift_reg48 (
        .clk           (clk),
        .rst_n         (rst_n),
        .shin_valid_i  (s48_shin_valid_i),
        .shin_data_i   (s48_shin_data_i),
        .sho_valid_o   (s48_sho_valid_o),
        .sho_data_o    (s48_sho_data_o)
    );

    assign s48_shin_valid_i = shin_valid_i;
    assign s48_shin_data_i = shin_data_i[(`SARRAY_LOAD_WIDTH/`SARRAY_H*49)-1:(`SARRAY_LOAD_WIDTH/`SARRAY_H*48)];
    assign sho_valid_o[48] = s48_sho_valid_o;
    assign sho_data_o[(`SARRAY_LOAD_WIDTH/`SARRAY_H*49)-1:(`SARRAY_LOAD_WIDTH/`SARRAY_H*48)] = s48_sho_data_o;



    // -------- shift_reg49

    wire [0:0]                                   s49_shin_valid_i;
    wire [`SARRAY_LOAD_WIDTH/`SARRAY_H-1:0]      s49_shin_data_i;
    wire [0:0]                                   s49_sho_valid_o;
    wire [`SARRAY_LOAD_WIDTH/`SARRAY_H-1:0]      s49_sho_data_o;

    shift_reg #(50) u_shift_reg49 (
        .clk           (clk),
        .rst_n         (rst_n),
        .shin_valid_i  (s49_shin_valid_i),
        .shin_data_i   (s49_shin_data_i),
        .sho_valid_o   (s49_sho_valid_o),
        .sho_data_o    (s49_sho_data_o)
    );

    assign s49_shin_valid_i = shin_valid_i;
    assign s49_shin_data_i = shin_data_i[(`SARRAY_LOAD_WIDTH/`SARRAY_H*50)-1:(`SARRAY_LOAD_WIDTH/`SARRAY_H*49)];
    assign sho_valid_o[49] = s49_sho_valid_o;
    assign sho_data_o[(`SARRAY_LOAD_WIDTH/`SARRAY_H*50)-1:(`SARRAY_LOAD_WIDTH/`SARRAY_H*49)] = s49_sho_data_o;



    // -------- shift_reg50

    wire [0:0]                                   s50_shin_valid_i;
    wire [`SARRAY_LOAD_WIDTH/`SARRAY_H-1:0]      s50_shin_data_i;
    wire [0:0]                                   s50_sho_valid_o;
    wire [`SARRAY_LOAD_WIDTH/`SARRAY_H-1:0]      s50_sho_data_o;

    shift_reg #(51) u_shift_reg50 (
        .clk           (clk),
        .rst_n         (rst_n),
        .shin_valid_i  (s50_shin_valid_i),
        .shin_data_i   (s50_shin_data_i),
        .sho_valid_o   (s50_sho_valid_o),
        .sho_data_o    (s50_sho_data_o)
    );

    assign s50_shin_valid_i = shin_valid_i;
    assign s50_shin_data_i = shin_data_i[(`SARRAY_LOAD_WIDTH/`SARRAY_H*51)-1:(`SARRAY_LOAD_WIDTH/`SARRAY_H*50)];
    assign sho_valid_o[50] = s50_sho_valid_o;
    assign sho_data_o[(`SARRAY_LOAD_WIDTH/`SARRAY_H*51)-1:(`SARRAY_LOAD_WIDTH/`SARRAY_H*50)] = s50_sho_data_o;



    // -------- shift_reg51

    wire [0:0]                                   s51_shin_valid_i;
    wire [`SARRAY_LOAD_WIDTH/`SARRAY_H-1:0]      s51_shin_data_i;
    wire [0:0]                                   s51_sho_valid_o;
    wire [`SARRAY_LOAD_WIDTH/`SARRAY_H-1:0]      s51_sho_data_o;

    shift_reg #(52) u_shift_reg51 (
        .clk           (clk),
        .rst_n         (rst_n),
        .shin_valid_i  (s51_shin_valid_i),
        .shin_data_i   (s51_shin_data_i),
        .sho_valid_o   (s51_sho_valid_o),
        .sho_data_o    (s51_sho_data_o)
    );

    assign s51_shin_valid_i = shin_valid_i;
    assign s51_shin_data_i = shin_data_i[(`SARRAY_LOAD_WIDTH/`SARRAY_H*52)-1:(`SARRAY_LOAD_WIDTH/`SARRAY_H*51)];
    assign sho_valid_o[51] = s51_sho_valid_o;
    assign sho_data_o[(`SARRAY_LOAD_WIDTH/`SARRAY_H*52)-1:(`SARRAY_LOAD_WIDTH/`SARRAY_H*51)] = s51_sho_data_o;



    // -------- shift_reg52

    wire [0:0]                                   s52_shin_valid_i;
    wire [`SARRAY_LOAD_WIDTH/`SARRAY_H-1:0]      s52_shin_data_i;
    wire [0:0]                                   s52_sho_valid_o;
    wire [`SARRAY_LOAD_WIDTH/`SARRAY_H-1:0]      s52_sho_data_o;

    shift_reg #(53) u_shift_reg52 (
        .clk           (clk),
        .rst_n         (rst_n),
        .shin_valid_i  (s52_shin_valid_i),
        .shin_data_i   (s52_shin_data_i),
        .sho_valid_o   (s52_sho_valid_o),
        .sho_data_o    (s52_sho_data_o)
    );

    assign s52_shin_valid_i = shin_valid_i;
    assign s52_shin_data_i = shin_data_i[(`SARRAY_LOAD_WIDTH/`SARRAY_H*53)-1:(`SARRAY_LOAD_WIDTH/`SARRAY_H*52)];
    assign sho_valid_o[52] = s52_sho_valid_o;
    assign sho_data_o[(`SARRAY_LOAD_WIDTH/`SARRAY_H*53)-1:(`SARRAY_LOAD_WIDTH/`SARRAY_H*52)] = s52_sho_data_o;



    // -------- shift_reg53

    wire [0:0]                                   s53_shin_valid_i;
    wire [`SARRAY_LOAD_WIDTH/`SARRAY_H-1:0]      s53_shin_data_i;
    wire [0:0]                                   s53_sho_valid_o;
    wire [`SARRAY_LOAD_WIDTH/`SARRAY_H-1:0]      s53_sho_data_o;

    shift_reg #(54) u_shift_reg53 (
        .clk           (clk),
        .rst_n         (rst_n),
        .shin_valid_i  (s53_shin_valid_i),
        .shin_data_i   (s53_shin_data_i),
        .sho_valid_o   (s53_sho_valid_o),
        .sho_data_o    (s53_sho_data_o)
    );

    assign s53_shin_valid_i = shin_valid_i;
    assign s53_shin_data_i = shin_data_i[(`SARRAY_LOAD_WIDTH/`SARRAY_H*54)-1:(`SARRAY_LOAD_WIDTH/`SARRAY_H*53)];
    assign sho_valid_o[53] = s53_sho_valid_o;
    assign sho_data_o[(`SARRAY_LOAD_WIDTH/`SARRAY_H*54)-1:(`SARRAY_LOAD_WIDTH/`SARRAY_H*53)] = s53_sho_data_o;



    // -------- shift_reg54

    wire [0:0]                                   s54_shin_valid_i;
    wire [`SARRAY_LOAD_WIDTH/`SARRAY_H-1:0]      s54_shin_data_i;
    wire [0:0]                                   s54_sho_valid_o;
    wire [`SARRAY_LOAD_WIDTH/`SARRAY_H-1:0]      s54_sho_data_o;

    shift_reg #(55) u_shift_reg54 (
        .clk           (clk),
        .rst_n         (rst_n),
        .shin_valid_i  (s54_shin_valid_i),
        .shin_data_i   (s54_shin_data_i),
        .sho_valid_o   (s54_sho_valid_o),
        .sho_data_o    (s54_sho_data_o)
    );

    assign s54_shin_valid_i = shin_valid_i;
    assign s54_shin_data_i = shin_data_i[(`SARRAY_LOAD_WIDTH/`SARRAY_H*55)-1:(`SARRAY_LOAD_WIDTH/`SARRAY_H*54)];
    assign sho_valid_o[54] = s54_sho_valid_o;
    assign sho_data_o[(`SARRAY_LOAD_WIDTH/`SARRAY_H*55)-1:(`SARRAY_LOAD_WIDTH/`SARRAY_H*54)] = s54_sho_data_o;



    // -------- shift_reg55

    wire [0:0]                                   s55_shin_valid_i;
    wire [`SARRAY_LOAD_WIDTH/`SARRAY_H-1:0]      s55_shin_data_i;
    wire [0:0]                                   s55_sho_valid_o;
    wire [`SARRAY_LOAD_WIDTH/`SARRAY_H-1:0]      s55_sho_data_o;

    shift_reg #(56) u_shift_reg55 (
        .clk           (clk),
        .rst_n         (rst_n),
        .shin_valid_i  (s55_shin_valid_i),
        .shin_data_i   (s55_shin_data_i),
        .sho_valid_o   (s55_sho_valid_o),
        .sho_data_o    (s55_sho_data_o)
    );

    assign s55_shin_valid_i = shin_valid_i;
    assign s55_shin_data_i = shin_data_i[(`SARRAY_LOAD_WIDTH/`SARRAY_H*56)-1:(`SARRAY_LOAD_WIDTH/`SARRAY_H*55)];
    assign sho_valid_o[55] = s55_sho_valid_o;
    assign sho_data_o[(`SARRAY_LOAD_WIDTH/`SARRAY_H*56)-1:(`SARRAY_LOAD_WIDTH/`SARRAY_H*55)] = s55_sho_data_o;



    // -------- shift_reg56

    wire [0:0]                                   s56_shin_valid_i;
    wire [`SARRAY_LOAD_WIDTH/`SARRAY_H-1:0]      s56_shin_data_i;
    wire [0:0]                                   s56_sho_valid_o;
    wire [`SARRAY_LOAD_WIDTH/`SARRAY_H-1:0]      s56_sho_data_o;

    shift_reg #(57) u_shift_reg56 (
        .clk           (clk),
        .rst_n         (rst_n),
        .shin_valid_i  (s56_shin_valid_i),
        .shin_data_i   (s56_shin_data_i),
        .sho_valid_o   (s56_sho_valid_o),
        .sho_data_o    (s56_sho_data_o)
    );

    assign s56_shin_valid_i = shin_valid_i;
    assign s56_shin_data_i = shin_data_i[(`SARRAY_LOAD_WIDTH/`SARRAY_H*57)-1:(`SARRAY_LOAD_WIDTH/`SARRAY_H*56)];
    assign sho_valid_o[56] = s56_sho_valid_o;
    assign sho_data_o[(`SARRAY_LOAD_WIDTH/`SARRAY_H*57)-1:(`SARRAY_LOAD_WIDTH/`SARRAY_H*56)] = s56_sho_data_o;



    // -------- shift_reg57

    wire [0:0]                                   s57_shin_valid_i;
    wire [`SARRAY_LOAD_WIDTH/`SARRAY_H-1:0]      s57_shin_data_i;
    wire [0:0]                                   s57_sho_valid_o;
    wire [`SARRAY_LOAD_WIDTH/`SARRAY_H-1:0]      s57_sho_data_o;

    shift_reg #(58) u_shift_reg57 (
        .clk           (clk),
        .rst_n         (rst_n),
        .shin_valid_i  (s57_shin_valid_i),
        .shin_data_i   (s57_shin_data_i),
        .sho_valid_o   (s57_sho_valid_o),
        .sho_data_o    (s57_sho_data_o)
    );

    assign s57_shin_valid_i = shin_valid_i;
    assign s57_shin_data_i = shin_data_i[(`SARRAY_LOAD_WIDTH/`SARRAY_H*58)-1:(`SARRAY_LOAD_WIDTH/`SARRAY_H*57)];
    assign sho_valid_o[57] = s57_sho_valid_o;
    assign sho_data_o[(`SARRAY_LOAD_WIDTH/`SARRAY_H*58)-1:(`SARRAY_LOAD_WIDTH/`SARRAY_H*57)] = s57_sho_data_o;



    // -------- shift_reg58

    wire [0:0]                                   s58_shin_valid_i;
    wire [`SARRAY_LOAD_WIDTH/`SARRAY_H-1:0]      s58_shin_data_i;
    wire [0:0]                                   s58_sho_valid_o;
    wire [`SARRAY_LOAD_WIDTH/`SARRAY_H-1:0]      s58_sho_data_o;

    shift_reg #(59) u_shift_reg58 (
        .clk           (clk),
        .rst_n         (rst_n),
        .shin_valid_i  (s58_shin_valid_i),
        .shin_data_i   (s58_shin_data_i),
        .sho_valid_o   (s58_sho_valid_o),
        .sho_data_o    (s58_sho_data_o)
    );

    assign s58_shin_valid_i = shin_valid_i;
    assign s58_shin_data_i = shin_data_i[(`SARRAY_LOAD_WIDTH/`SARRAY_H*59)-1:(`SARRAY_LOAD_WIDTH/`SARRAY_H*58)];
    assign sho_valid_o[58] = s58_sho_valid_o;
    assign sho_data_o[(`SARRAY_LOAD_WIDTH/`SARRAY_H*59)-1:(`SARRAY_LOAD_WIDTH/`SARRAY_H*58)] = s58_sho_data_o;



    // -------- shift_reg59

    wire [0:0]                                   s59_shin_valid_i;
    wire [`SARRAY_LOAD_WIDTH/`SARRAY_H-1:0]      s59_shin_data_i;
    wire [0:0]                                   s59_sho_valid_o;
    wire [`SARRAY_LOAD_WIDTH/`SARRAY_H-1:0]      s59_sho_data_o;

    shift_reg #(60) u_shift_reg59 (
        .clk           (clk),
        .rst_n         (rst_n),
        .shin_valid_i  (s59_shin_valid_i),
        .shin_data_i   (s59_shin_data_i),
        .sho_valid_o   (s59_sho_valid_o),
        .sho_data_o    (s59_sho_data_o)
    );

    assign s59_shin_valid_i = shin_valid_i;
    assign s59_shin_data_i = shin_data_i[(`SARRAY_LOAD_WIDTH/`SARRAY_H*60)-1:(`SARRAY_LOAD_WIDTH/`SARRAY_H*59)];
    assign sho_valid_o[59] = s59_sho_valid_o;
    assign sho_data_o[(`SARRAY_LOAD_WIDTH/`SARRAY_H*60)-1:(`SARRAY_LOAD_WIDTH/`SARRAY_H*59)] = s59_sho_data_o;



    // -------- shift_reg60

    wire [0:0]                                   s60_shin_valid_i;
    wire [`SARRAY_LOAD_WIDTH/`SARRAY_H-1:0]      s60_shin_data_i;
    wire [0:0]                                   s60_sho_valid_o;
    wire [`SARRAY_LOAD_WIDTH/`SARRAY_H-1:0]      s60_sho_data_o;

    shift_reg #(61) u_shift_reg60 (
        .clk           (clk),
        .rst_n         (rst_n),
        .shin_valid_i  (s60_shin_valid_i),
        .shin_data_i   (s60_shin_data_i),
        .sho_valid_o   (s60_sho_valid_o),
        .sho_data_o    (s60_sho_data_o)
    );

    assign s60_shin_valid_i = shin_valid_i;
    assign s60_shin_data_i = shin_data_i[(`SARRAY_LOAD_WIDTH/`SARRAY_H*61)-1:(`SARRAY_LOAD_WIDTH/`SARRAY_H*60)];
    assign sho_valid_o[60] = s60_sho_valid_o;
    assign sho_data_o[(`SARRAY_LOAD_WIDTH/`SARRAY_H*61)-1:(`SARRAY_LOAD_WIDTH/`SARRAY_H*60)] = s60_sho_data_o;



    // -------- shift_reg61

    wire [0:0]                                   s61_shin_valid_i;
    wire [`SARRAY_LOAD_WIDTH/`SARRAY_H-1:0]      s61_shin_data_i;
    wire [0:0]                                   s61_sho_valid_o;
    wire [`SARRAY_LOAD_WIDTH/`SARRAY_H-1:0]      s61_sho_data_o;

    shift_reg #(62) u_shift_reg61 (
        .clk           (clk),
        .rst_n         (rst_n),
        .shin_valid_i  (s61_shin_valid_i),
        .shin_data_i   (s61_shin_data_i),
        .sho_valid_o   (s61_sho_valid_o),
        .sho_data_o    (s61_sho_data_o)
    );

    assign s61_shin_valid_i = shin_valid_i;
    assign s61_shin_data_i = shin_data_i[(`SARRAY_LOAD_WIDTH/`SARRAY_H*62)-1:(`SARRAY_LOAD_WIDTH/`SARRAY_H*61)];
    assign sho_valid_o[61] = s61_sho_valid_o;
    assign sho_data_o[(`SARRAY_LOAD_WIDTH/`SARRAY_H*62)-1:(`SARRAY_LOAD_WIDTH/`SARRAY_H*61)] = s61_sho_data_o;



    // -------- shift_reg62

    wire [0:0]                                   s62_shin_valid_i;
    wire [`SARRAY_LOAD_WIDTH/`SARRAY_H-1:0]      s62_shin_data_i;
    wire [0:0]                                   s62_sho_valid_o;
    wire [`SARRAY_LOAD_WIDTH/`SARRAY_H-1:0]      s62_sho_data_o;

    shift_reg #(63) u_shift_reg62 (
        .clk           (clk),
        .rst_n         (rst_n),
        .shin_valid_i  (s62_shin_valid_i),
        .shin_data_i   (s62_shin_data_i),
        .sho_valid_o   (s62_sho_valid_o),
        .sho_data_o    (s62_sho_data_o)
    );

    assign s62_shin_valid_i = shin_valid_i;
    assign s62_shin_data_i = shin_data_i[(`SARRAY_LOAD_WIDTH/`SARRAY_H*63)-1:(`SARRAY_LOAD_WIDTH/`SARRAY_H*62)];
    assign sho_valid_o[62] = s62_sho_valid_o;
    assign sho_data_o[(`SARRAY_LOAD_WIDTH/`SARRAY_H*63)-1:(`SARRAY_LOAD_WIDTH/`SARRAY_H*62)] = s62_sho_data_o;



    // -------- shift_reg63

    wire [0:0]                                   s63_shin_valid_i;
    wire [`SARRAY_LOAD_WIDTH/`SARRAY_H-1:0]      s63_shin_data_i;
    wire [0:0]                                   s63_sho_valid_o;
    wire [`SARRAY_LOAD_WIDTH/`SARRAY_H-1:0]      s63_sho_data_o;

    shift_reg #(64) u_shift_reg63 (
        .clk           (clk),
        .rst_n         (rst_n),
        .shin_valid_i  (s63_shin_valid_i),
        .shin_data_i   (s63_shin_data_i),
        .sho_valid_o   (s63_sho_valid_o),
        .sho_data_o    (s63_sho_data_o)
    );

    assign s63_shin_valid_i = shin_valid_i;
    assign s63_shin_data_i = shin_data_i[(`SARRAY_LOAD_WIDTH/`SARRAY_H*64)-1:(`SARRAY_LOAD_WIDTH/`SARRAY_H*63)];
    assign sho_valid_o[63] = s63_sho_valid_o;
    assign sho_data_o[(`SARRAY_LOAD_WIDTH/`SARRAY_H*64)-1:(`SARRAY_LOAD_WIDTH/`SARRAY_H*63)] = s63_sho_data_o;



endmodule