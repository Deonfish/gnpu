module shift_reg(
	input 							 clk,
	input 							 rst_n,
	input  [0:0] 					 shin_valid_i,
	input  [`SARRAY_LOAD_WIDTH-1:0]  shin_data_i,
	output [`SARRAY_H-1:0] 			 sho_valid_o,
	output [``SARRAY_LOAD_WIDTH-1:0] sho_data_o
);


endmodule